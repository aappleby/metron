module Module
(
);
/*public:*/
endmodule
