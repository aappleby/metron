`include "metron_tools.sv"

