`ifndef METRON_H_SV
`define METRON_H_SV

/* verilator lint_off width */
/* verilator lint_off IGNOREDRETURN */

`default_nettype none

typedef int unsigned uint32_t;
typedef int int32_t;

`endif
