`include "metron/metron_tools.sv"

// We need to support very basic preprocessor macros or else dealing with mixed
// languages will be a huge pain in the butt.

#ifdef METRON_SV

//module Submod();
//endmodule

#else

`endif

/*
#endif


#ifndef METRON_SV

#else

#endif


#ifdef METRON_CPP

#else

#endif
*/
