`include "metron/tools/metron_tools.sv"

module Module (
{{port list}}
);
/*public:*/

  LSKJLKDJF
{{13CNodeFunction}}

  {{13CNodeFunction}}

/*private:*/

  logic x;
  logic y;
  logic z;
  logic[1:0] out;
endmodule;