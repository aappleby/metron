`include "metron/tools/metron_tools.sv"
