// This file should always fail in everything

module Module (input logic clock);
  always_ff @ (posedge clock) begin
    af8902h[f0a9sdj'[pfjioa'sdjfalsdknvzx,.cmnvz/xvjk"v0[p2qui]30-9fa]09sdiuf'sj
  end
endmodule
