`include "metron_tools.sv"

// Empty module should pass.

module Module
(
input logic clock
);

endmodule
