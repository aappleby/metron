`include "metron/tools/metron_tools.sv"

// Empty module should pass.

module Module  (
);
endmodule
