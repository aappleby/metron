`include "metron_tools.sv"

// Getter methods should turn into outputs.

module Module
(
  input logic clock,
  output logic[6:0] get_reg_ret
);
/*public:*/

  function logic[6:0] get_reg();
    get_reg = my_reg;
  endfunction
  always_comb get_reg_ret = get_reg();

  always_comb begin : tock
  end


/*private:*/

  task automatic tick();
    my_reg <= my_reg + 1;
  endtask
  always_ff @(posedge clock) tick();

  logic[6:0] my_reg;
endmodule
