// Comments at start of file should be preserved

`include "metron/tools/metron_tools.sv"

// Empty module should pass.

module Module (
);
endmodule

// Comments at end of file should be preserved
