`include "metron_tools.sv"

module Module
(
input logic clock
);
endmodule

