`include "metron_tools.sv"

// Increment/decrement should _not_ return a value.

module Module
(
input logic clock
);
/*public:*/
endmodule

