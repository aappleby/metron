`include "metron/tools/metron_tools.sv"

module Module (
);
/*public*/

  parameter q = 7;
  initial begin
    x = 1;
    y = 2;
    z = 3;
  end

/*private*/

  /*logic<1> x;*/
  /*logic<1> y;*/
  /*logic<1> z;*/
  /*logic<2> out;*/
endmodule
