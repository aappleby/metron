module Top (
{{port list}}
);
{{template parameter list}}
/*public:*/
endmodule;