`include "metron/metron_tools.sv"
