`include "metron_tools.sv"

// Namespaces turn into packages.
// "using" doesn't work in methods right now :/

package MyPackage;
  parameter int foo = 3;
endpackage

module Module
(
  input logic clock,
  output int my_sig,
  output int my_reg,
  output int tock_ret
);
/*public:*/


  always_comb begin : tock
    my_sig = MyPackage::foo + 1;
    tock_ret = my_sig;
  end

  task automatic tick();
    my_reg <= my_reg + MyPackage::foo;
  endtask
  always_ff @(posedge clock) tick();
endmodule
