`include "metron_tools.sv"

module Pong
(
	input logic clock
);
/*public:*/

	always_comb begin /*tock*/
	end

/*private:*/
endmodule




